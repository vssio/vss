module paths

import net.urllib

fn add_context_root(base_url string, relative_path string) string {
	return ''
}
